module digital_clock_top_tb();
    reg        clk;
    reg        rst_n;
    reg  [6:0] key;
    
    wire [5:0] sel;                   //数码管位选（选择当前要显示的数码管）
	wire [6:0] seg;                   //数码管段选（当前要显示的内容） 
    wire       time_led;
    wire       beep;
    
    //---- key0 日期，时间切换
    //---- key1 模式切换 （时钟，闹钟，秒表，调时）
    //---- key2 调时和设置闹钟时，小时、分钟左右切捯
    //---- key3 +1 
    //---- key4 -1
    //---- key5 秒表暂停（开始）切换
    //---- key6 秒表清除
    
    initial clk = 0;
    always #1 clk = ~clk;
    
    initial begin
        rst_n = 0;
        key = 7'b1111111;
        #10;
        key[0] = 0;   // 显示日期
        #30;           // 按键低电平持续一段时间，防止被filter滤掉
        key[0] = 1;
        #100;
        key[0] = 0;  // 正常显示时间
        #30;       
        key[0] = 1;
//------------------------------------------ 设置闹钟 -------------------------------------------------------
        #1000;
        key[1] = 0;    //闹钟模式
        #30;       
        key[1] = 1;
        #5;
        
        repeat(20) begin  //分个位+
            #20;
            key[3] = 0; 
            #30;       
            key[3] = 1;    
        end
        
        #5;
        key[2] = 0;      //分十位
        #30;       
        key[2] = 1;
        repeat(12) begin  //分十位+
            #20;
            key[3] = 0; 
            #30;       
            key[3] = 1;    
        end
        
        #5;
        key[2] = 0;      //小时个位
        #30;       
        key[2] = 1;
        repeat(24) begin  //小时个位+   
            #20;
            key[3] = 0; 
            #30;       
            key[3] = 1;    
        end 
     // 闹钟设置为24:00:00
//------------------------------------------ 秒表模式 -------------------------------------------------------
        #1000;
        key[1] = 0;    //秒表模式
        #30;       
        key[1] = 1;
        #5;
        
        key[5] = 0;   //开始  
        #30;       
        key[5] = 1;
        #5;
        
        key[5] = 0;   //暂停  
        #30;       
        key[5] = 1;
        #5;
        
        key[5] = 0;   //开始  
        #30;       
        key[5] = 1;
        #5;
        
        key[6] = 0;   //清除  
        #30;       
        key[6] = 1;
        #5;
//------------------------------------------ 校准时间 -------------------------------------------------------        
        #5;
        key[1] = 0;  
        #30;       
        key[1] = 1;
        #5;
        
        repeat(61) begin  //校准秒位+
            #20;
            key[3] = 0; 
            #30;       
            key[3] = 1;    
        end
        repeat(61) begin  //校准秒位-
            #20;
            key[4] = 0; 
            #30;       
            key[4] = 1;    
        end
        
        #10;
        key[2] = 0;    //校准分位
        #30;       
        key[2] = 1;
        
        repeat(61) begin  //校准分位+
            #20;
            key[3] = 0; 
            #30;       
            key[3] = 1;    
        end
        repeat(61) begin  //校准分位-
            #20;
            key[4] = 0; 
            #30;       
            key[4] = 1;    
        end
        
        #10;
        key[2] = 0;    //校准小时位
        #30;       
        key[2] = 1;
        
        repeat(61) begin  //校准小时位+
            #20;
            key[3] = 0; 
            #30;       
            key[3] = 1;    
        end
        repeat(61) begin  //校准小时位-
            #20;
            key[4] = 0; 
            #30;       
            key[4] = 1;    
        end
        
        
        
        
        
    end
    
    digital_clock_top UU1(
            .clk            (clk),
            .rst_n          (rst_n),
            .key_in         (key),
            .sel            (sel), 
            .seg            (seg),   
            .time_led       (time_led),
            .beep           (beep)
    );

endmodule